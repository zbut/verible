// 'localparams' should only be declared within modules' and classes' definition bodies.
// verilog_lint: waive parameter-name-prefix
localparam int Foo = 1;
