// Expect the parameter to explicitly define a storage type
// verilog_lint: waive parameter_name_prefix
parameter Bar = 1;
