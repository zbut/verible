// Expected parameter name, "Hello_World" to follow UpperCamelCase or ALL_CAPS naming convention.
// verilog_lint: waive parameter_name_prefix
parameter int Hello_World = 1;
