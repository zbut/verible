parameter int HELLO_WORLD = 1;
