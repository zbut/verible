// Expect the parameter to explicitly define a storage type
// verilog_lint: waive parameter-name-prefix
parameter Bar = 1;
