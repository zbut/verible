// Expected parameter type name, "Hello_World" to follow lower_snake_case naming convention and end with _t.
// verilog_lint: waive parameter-name-prefix
parameter type Hello_World = logic;
