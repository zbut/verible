// 'localparams' should only be declared within modules' and classes' definition bodies.
// verilog_lint: waive parameter-name-prefix
// verilog_lint: waive parameter-name-style
localparam int Foo = 1;
