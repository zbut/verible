parameter int P_HELLO_WORLD = 1;
