// Expect the parameter to explicitly define a storage type
// verilog_lint: waive parameter-name-prefix
// verilog_lint: waive parameter-name-style
parameter Bar = 1;
