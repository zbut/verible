// 'localparams' should only be declared within modules' and classes' definition bodies.
// verilog_lint: waive parameter_name_prefix
localparam int Foo = 1;
