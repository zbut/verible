module port_name_style(input bit hello_world_i);
endmodule
